module top_module ( input a, input b, output out );

    mod_a mod_a_obj(a, b, out);
    
endmodule
